
typedef strcut packed{
   logic [10:0] bits;
   } encoder_t

typedef strcut packed{
   logic [11:0] bits;
   } decoder_t  
